-- -----------------------------------------------------------------
-- "Copyright (C) Altium Limited 2003"
-- -----------------------------------------------------------------
-- Component Name: 	BUFE16B
-- Description: 	16-Bit 3-state Buffer with Active High Enable, Bus Version
-- Core Revision: 	1.00.00
-- -----------------------------------------------------------------
-- Modifications with respect to Version  : 
--
--
-- -----------------------------------------------------------------

LIBRARY ieee;
    USE ieee.std_logic_1164.ALL;

-- -----------------------------------------------------------------
-- Entity for BUFE16B
-- -----------------------------------------------------------------
ENTITY BUFE16B IS
    Port(	E: IN std_logic:='U';
    		I: IN  std_logic_vector(15 downto 0):=(others => 'U');
         	O: OUT std_logic_vector(15 downto 0));
end BUFE16B;
-- -----------------------------------------------------------------

-- -----------------------------------------------------------------
-- Architecture behav for BUFE16B
-- -----------------------------------------------------------------
ARCHITECTURE behav OF BUFE16B IS
-- -----------------------------------------------------------------
-- -----------------------------------------------------------------
begin
-- -----------------------------------------------------------------

   O <= I when E='1' else (others => 'Z');
-- -----------------------------------------------------------------
end behav;
-- -----------------------------------------------------------------
